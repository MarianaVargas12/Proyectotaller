module condcheck();

endmodule 