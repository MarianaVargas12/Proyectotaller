module condlogic();

endmodule 